
module myhardware (
	reset_reset_n,
	clk_clk,
	leds_export,
	hex0_export,
	hex1_export,
	hex2_export,
	hex3_export,
	hex4_export,
	hex5_export);	

	input		reset_reset_n;
	input		clk_clk;
	output	[9:0]	leds_export;
	output	[6:0]	hex0_export;
	output	[6:0]	hex1_export;
	output	[6:0]	hex2_export;
	output	[6:0]	hex3_export;
	output	[6:0]	hex4_export;
	output	[6:0]	hex5_export;
endmodule
